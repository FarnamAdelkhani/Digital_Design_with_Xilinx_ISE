-- Vhdl test bench created from schematic C:\Users\User_Account\Desktop\test\Lab7\labo7part3.sch - Tue Mar 03 15:41:31 2015
--
-- Notes: 
-- 1) This testbench template has been automatically generated using types
-- std_logic and std_logic_vector for the ports of the unit under test.
-- Xilinx recommends that these types always be used for the top-level
-- I/O of a design in order to guarantee that the testbench will bind
-- correctly to the timing (post-route) simulation model.
-- 2) To use this template as your testbench, change the filename to any
-- name of your choice with the extension .vhd, and use the "Source->Add"
-- menu in Project Navigator to import the testbench. Then
-- edit the user defined section below, adding code to generate the 
-- stimulus for your design.
--
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
LIBRARY UNISIM;
USE UNISIM.Vcomponents.ALL;
ENTITY labo7part3_labo7part3_sch_tb IS
END labo7part3_labo7part3_sch_tb;
ARCHITECTURE behavioral OF labo7part3_labo7part3_sch_tb IS 

   COMPONENT labo7part3
   PORT( );
   END COMPONENT;


BEGIN

   UUT: labo7part3 PORT MAP(
		
   );

-- *** Test Bench - User Defined Section ***
   tb : PROCESS
   BEGIN
      WAIT; -- will wait forever
   END PROCESS;
-- *** End Test Bench - User Defined Section ***

END;
